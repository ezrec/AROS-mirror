En bunt AROS-utvecklare och AROS-fans, i ett soligt och väldigt hett Naples.
