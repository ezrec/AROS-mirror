På semester i Djerba, Tunisien
