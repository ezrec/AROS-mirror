=============
Status Update
=============

:Author:   Paolo Besser
:Date:     2007-10-01

Senaste nyheter
---------------

Nyhet! Neil Cafferkey har bidragit med en helt ny `installer`__ f�r
AROS, vilket m�jligg�r en renare och s�krare installation p� h�rddiskar.
Nya finnesser enligt nedan:

- Installationsdisk och partitioner kan nu anges.
- Skapandet av en Work-partition fungerar.
- Partitionsstorlekar kan anges och existerande partitioner kan beh�llas.
- Windows �r tillagd till GRUB boot menu om en existerande Windows-partition hittas.


Notera dock, att detta fortfarande �r en beta-version. H�r f�ljer n�gra
varningar fr�n Neil: " Den nya h�rddisk-installern �r nu inkluderad
i "Nightly ISO" och �r f�rdig f�r testning. Men, det finns f�r tillf�llet
en bug i antingen Wanderer eller FFS som m�ste �tg�rdas. Efter att man startat
installern, s� m�ste du avsluta Wanderer innan du forts�tter (om du inte
kommer att formatera n�gon partition).
Var extra f�rsiktig �n vanligt med denna version av installern, uts�tt inte
datorn med ej s�kerhetskopierad data. Den borde beh�lla alla existerande
partitioner, men inte s� m�nga har testat detta f�rutom jag."

Om du har en testdator med ej viktig data p�, s� vore det b�sta om du
laddar ner 10-01 "nightly build (eller senare) och hj�lper oss att hitta
buggar. Du kan anv�nda Bug Tracker eller skicka ett meddelande i detta
AROS-Exec `discussion`__. 

Demonstration av AROS
---------------------

Som tidigare n�mnt p� denna hemsida s� har AROS varit en g�ststj�rna p�
`Pianeta Amiga 2007`__.  Under den popul�ra amigashowen s� har
Paulo Besser presenterat AROS till en del intresserade Amiga-anh�ngare.
Evenemanget har n�mnts i n�gra st�rre IT-nyhets-hemsidor som `TGM Online`__
och `HW Upgrade`__. En rapport av evenemanget har blivit publicerad av 
`The AROS Show`__ (L�s denna `here`__) Du kan �ven se en trevlig `video`__
p� YouTube.

__ http://mama.indstate.edu/users/nova/installer.jpg
__ http://aros-exec.org/modules/newbb/viewtopic.php?topic_id=2319
__ http://www.pianetaamiga.it/2007/eng/
__ http://tgmonline.futuregamer.it/news/settembre2007/20070910111905
__ http://www.hwupgrade.it/news/videogiochi/presentazione-italiana-per-l-os-indipendente-aros_22619-0.html
__ http://arosshow.blogspot.com
__ http://arosshow.blogspot.com/2007/09/pianeta-amiga-2007-report-from-paolo.html
__ http://video.google.it/videoplay?docid=-3563710058663289244
