Tack vare Sergey Mineychev, så är alla AROS-programmens cataloger lokaliserade samt att typsnitten är inlagda (med tillstånd av Michael Malyshev, ATO).
