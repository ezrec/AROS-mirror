.. raw:: html

   <h1>Introduktion<br><img style="width: 238px; height: 2px;" alt="spacer" src="/images/sidespacer.png"></h1>

.. raw:: html

  <?php include('../rsfeed/randimg.php');  random_image("/images/thubs/","100","76"); ?>

AROS �r ett portabelt och fritt operativsystem f�r desktop med syfte p�
att vara kompatibelt med AmigaOS 3.1, och samtidigt f�rb�ttra det i
m�nga omr�den. K�llkoden �r tillg�nglig under en open source-licens, vilket
till�ter alla friheten att f�rb�ttra det.
