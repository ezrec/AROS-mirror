Michael Schultz arbetandes i MADIREL-laboratoriet i Marsiell/Frankrike med
någon typ av elektroder.
