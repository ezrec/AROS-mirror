Tack vare Michal Schultz så har AROS nu ett fungerande PCI-stöd. Denna skärmdump
visar PCITool, ett program som låter dig browsa i en lista av alla PCI-devices
som sitter i din dator.
