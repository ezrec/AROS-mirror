På tur i de norska fjällen.
