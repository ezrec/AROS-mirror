=================
Tillk�nnagivanden
=================

Denna produkt inneh�ller mjukvara utvecklad av University of California,
Berkeley och deras medarbetare.

Denna mjukvara �r delvis baserad p� arbeten fr�n the Independent JPEG Group.

Denna mjukvara �r delvis baserad p� arbeten fr�n the FreeType Team.

Denna mjukvara �r delvis baserad p� arbeten fr�n Catharon Productions, Inc.

Graphics Interchange Format(c) �r upphovsr�ttskyddad egendom tillh�rande CompuServer Incorporated.
GIF(sm) �r ett Service Mark tillh�rande CompuServer Incorporated.
