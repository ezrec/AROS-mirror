===========
Nerladdning
===========

.. Contents::

.. Note::

   När du laddar ner "nightly builds", så måste du använda en nerladdnings-
   hanterare så att du kan återuppta en avbruten nerladdning, eller en
   textbaserad applikation som t.ex. wget (Du kan använda "wget -c" för
   att återuppta nerladdningen av en fil som är nerladdad av ett annat program).

Snapshots
=========

Från den 1:a mars 2007 är snapshots av AROS inte längre tillgängliga. Vi
uppmanar alla som vill testa AROS att ladda ner den senaste "nightly build"
istället. AROS växer väldigt fort, och snapshots innehåller oftast
föråldad kod. Vi tror också att "nightly builds" är mer användbara med 
tanke på betatestningen: använd gärna `bug tracker`__ för att rapportera buggar.

__ http://sourceforge.net/tracker/?atid=439463&group_id=43586&func=browse


Nightly builds
==============

"Nightly builds" görs, som man ser på namnet, automatiskt varje natt direkt
från subversions-trädet och innehåller den senaste koden. Men dessa har inte
blivit testade och kan innehålla buggar. Dock fungerar dom för det mesta bra.

Rapportera gärna buggar som du hittar när du använder "nightly builds" till
`bug tracker`__. För övriga ärenden eller frågor, kontakta oss via
`AROS-Exec`__ forumen.

.. raw:: html

   <?php virtual( "/cgi-bin/files?type=nightly&lang=en" ); ?>

__ http://sourceforge.net/tracker/?atid=439463&group_id=43586&func=browse
__ http://aros-exec.org/

