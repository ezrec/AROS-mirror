Denna skärmdump visar den kommande GUI FTP-klienten av voidstar aka suppah, tagen från den senaste builden.
