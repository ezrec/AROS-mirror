P� semester i Djerba, Tunisien
