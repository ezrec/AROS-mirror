=================
Statusuppdatering
=================

:F�rfattare:   Paolo Besser
:Datum:     2006-08-28

Aros.org finns nu tillg�nglig i ytterligare tv� spr�k: tack vare Sergey Mineychew
kan du nu se hemsidan p� `Rysska`__, medans Tomasz Paul fortfarande jobbar p� den
`Polska`__ �vers�ttningen. Du beh�ver bara klicka i menyn i �vre v�nstra h�rnet
f�r att n� de nya sidorna. Sergey jobbar ocks� med Rysska locales till 
AROS-applikationer.

__ http://www.aros.org/ru/index.php
__ http://www.aros.org/pl/index.php

