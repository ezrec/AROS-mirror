Zune blir bara b�ttre och b�ttre! Nu tack vare Georg Steger s� har
vi fler classes implementerade, som du kan se. Du kan �ven se gcc
kompilera ett av test-programmen f�r de nya implementerade classes.
