
.. Include:: introduction/index-abstract.sv

`L�s mer... <introduction/index>`__

.. Include:: documentation/developers/contribute-abstract.sv

`L�s mer... <documentation/developers/contribute>`__

.. Include:: news/index.sv
