Mer sidor i Zune-inst�llningarna.
