Matt "Crazy" Parsons som observerar Hubble space teleskopet.
