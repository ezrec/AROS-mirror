===========
Skärmdumpar
===========

