H�r har vi n�gra nya funktioner i icon-library. Du kan se den nya effekten 
f�r de valda ikonerna ("S"-mappen �r vald h�r, d�rf�r �r den ljusare �n de
andra ikonerna). Ikon-namnen ritas nu upp med en outline, f�r att bli 
synliga �ven p� en m�rk bakgrund (detta kommer naturligtvis �ven att vara
konfigurerbart f�r anv�ndarna i framtiden).

Vi kan �ven se fil-identifikationen i bruk: text-filerna i "S"-mappen f�r
speciella def_Text-ikoner, medans filen "AROS.png" f�r den generella
projekt-ikonen. Vi har inte s� m�nga ikoner just nu, men om de fanns
tillg�ngliga s� skulle "AROS.png" f� en def_Picture-ikon (Eller �ven kanske
en def_PNG-ikon om det fanns tillg�ngligt).
