P� jobbet.
