Om du n�gonsin undrat �ver hur Fabias ansikte ser ut, s� vet du det nu! :)
