N�gra enkla demos av den tidiga (och i utveckling) Mesa-portningen.
