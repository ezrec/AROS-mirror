Denna sk�rmdump visar den kommande GUI FTP-klienten av voidstar aka suppah, tagen fr�n den senaste builden.
