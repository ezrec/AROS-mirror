Distributioner
==============

Distributioner �r konfigurerade och testade versioner av AROS.
Dom inneh�ller en m�ngd anv�ndarprogram som inte finns med i dom vanliga AROS.org utg�vorna. Dessa distributioner riktar sig till fr�mst till intresserade anv�ndare. Dessa har ev. inte dom senaste k�rn uppdateringarna, men anv�ndar v�nligheten och stabiliteten �r betydligt st�rre, �n f�r dom nattliga utg�vorna. 

Om du �r en anv�ndare som �r intresserad av AROS, s� rekomenderar vi att du b�rjar med den senaste distributionen, f�r att f� den b�sta m�jliga erfarenheten av AROS systemet.
