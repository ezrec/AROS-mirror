=================
Statusuppdatering
=================

:F�rfattare:   Paolo Besser
:Datum:     2006-06-20

Tack vare Matthias Rustlers s� finns aros.org nu ocks� p� `Tyska`__, vilken
du hittar p� www.aros.org/de/.
Men du beh�ver inte komma ih�g varje spr�ks hemsida eftersom
vi har lagt till en internationell meny p� v�nstersidan. Bara v�lj ditt
favoritspr�k och skapa ett bokm�rke f�r bekv�m �tkomst.

__ http://www.aros.org/de/index.php



New PPC snapshot!
-----------------

There is a new binary snapshot for hosted AROS-PPC! Just go to Sourceforge 
website and `download it`__! Here's the release notes: "This release depends 
on glibc 2.3.2 or newer. You need to give AROS some more RAM than the default 
allocation of 16 MB (leaves about 4 MB for applications). Start it using: 
./aros -m 64 This will allocate 64 MB. As with all X11 hosted AROS versions 
you need to add Option "BackingStore" to the Device section of xorg.conf"


__ http://sourceforge.net/project/shownotes.php?group_id=43586&release_id=425583
