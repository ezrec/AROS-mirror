Michael Schultz arbetandes i MADIREL-laboratoriet i Marsiell/Frankrike med
n�gon typ av elektroder.
