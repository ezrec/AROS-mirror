Väntar som många andra på Amiga Inc på WoA 1999.
