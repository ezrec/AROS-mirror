=================
Statusuppdatering
=================

:F�rfattare:   Paolo Besser
:Datum:     2006-09-15

�vers�ttningen av aros.org forts�tter. Samuel Atlan jobbar p� sin
`Franska �vers�ttning`__ av v�r hemsida. Det kommer att ta lite tid
innan det blir f�rdigt men de f�rsta sidorna finns redans tillg�ngliga
fr�n menyn i �vre v�nstra h�rnet. Nytt p� aros.org �r ocks� att man
nu kan n� de �versatta sidorna genom att l�gga till spr�kkoden efter 
den vanliga URL-en. Som exempel hittar du den Italienska sidan under
*www.aros.org/it*, den Ryska p� *www.aros.org/ru* och s� vidare.

__ http://www.aros.org/fr/

AROS i nyheterna
----------------

Vi rekommenderar den h�r trevliga `recensionen`__ som Dmitar Butrovski har
skrivit p� `OSnews.com`__. Det �r utan tvekan en av de mest kompletta artiklar
som har skrivits om v�rat fina operativsystem. Om du inte redan �r bekant med
vad AROS �r s� f�r du antagligen en bra id� om det.

__ http://osnews.com/story.php?news_id=15819
__ http://osnews.com

Mjukvara
--------

Version 1.20 av den *VICE*, den ber�mda emulatorn av Commodores linje av
8-bitars datorer, finns nu tillg�nglig f�r alla Amiga-plattformar inklusive AROS.
Du hittar den `h�r`__.

*WinAros* �r en f�rinstallerad AROS-milj� installerad p� en h�rddisk-avbildning,
kompatibel med de v�lk�nda virtualiseringsmilj�erna QEMU och Microsoft
VirtualPC, b�da fritt tillg�ngliga p� Internet. Du kan ladda ner 
`QEMU Winaros h�r`__ och `QEMU VirtualPC h�r`__. Heinz-Raphael Reinke har ocks�
skrivit en komplett guide �ver `AROS-installation p� h�rddisk`__ i PDF-format.
Den finns �ven p� `Tyska`__ om du f�redrar det. Du beh�ver Adobe Acrobat
Reader, FoxIt Reader eller aPDF/xPDF f�r att l�sa dem.

*Installation Kit for AROS (IKAROS)* �r en upps�ttning med h�rddisk-avbildningar
f�r olika virtualiseringsmilj�er, s�som QEMU och VMWare, redan partitionerade,
formatterade och f�rdiga att installera AROS p�. F�rdelarna med det �r liten 
storlek p� arkiven man laddar hem eftersom den inte beh�ver stora m�ngder med filer,
och m�jligheten att installera nya, fr�sha versioner av AROS. Det g�r det enkelt
att testa nattliga kompileringar utan att beh�va st�ka med partitionering.
Instruktioner �ver hur man installerar medf�ljer.
V�nligen bes�k `Aros-Exec`__ f�r uppdateringar och nerladdning.

__ http://www.viceteam.org/amigaos.html
__ http://amidevcpp.amiga-world.de/WinAros/WinAros_Light_QEMU.zip
__ http://amidevcpp.amiga-world.de/WinAros/WinAros_Light_VPC.zip
__ http://amidevcpp.amiga-world.de/WinAros/Aros_HD_Install_English.pdf
__ http://amidevcpp.amiga-world.de/WinAros/Aros_HD_Installation.pdf
__ http://archives.aros-exec.org/?function=showfile&file=emulation/misc/arosik02.zip
