========
L�nkning
========

:Author:    Adam Chodorowski
:Copyright: Copyright � 2001-2007, The AROS Development Team
:Version:   $Revision$
:Date:      $Date$
:Status:    Done.

Ett mycket bra s�tt att visa ditt st�d f�r AROS, och f�r att uppmana andra,
�r att l�nka till denna hemsida fr�n din egen. Du kan anv�nda en av nedanst�ende banners
f�r detta �ndam�l.

+------------------------------------------+----------------------+
| Bild                                     | Upphovsman           |
+==========================================+======================+
| .. Image:: /images/aros-banner.gif       | Cyb0rg / Resistance  |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-banner2.png      | S33k_100             |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-banner-blue.png  | S33k_100             |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-banner-pb2.png   | Paolo Besser         |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-banner-peta.png  | Petr Novak           |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+


Alternativt s� finns det �ven signatur-banners f�r anv�ndning i forum:

+------------------------------------------+----------------------+
| Bild                                     | Upphovsman           |
+==========================================+======================+
| .. Image:: /images/aros-sigbar-user.png  | S33k_100             |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-sigbar-coder.png | S33k_100             |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+


Var v�nlig, l�nka direkt till http://www.aros.org/ och inte till n�gon av de speglade
hemsidorna eftersom dessa kan �ndras. Se �ven till att ha en lokal kopia av bilden f�r
att minska bandbredden.
