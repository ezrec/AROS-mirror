P� tur i de norska fj�llen.
