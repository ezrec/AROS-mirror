===========
Sk�rmdumpar
===========

