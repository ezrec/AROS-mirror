Tack vare Michal Schultz s� har AROS nu ett fungerande PCI-st�d. Denna sk�rmdump
visar PCITool, ett program som l�ter dig browsa i en lista av alla PCI-devices
som sitter i din dator.
