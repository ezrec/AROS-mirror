Vi beh�ver din hj�lp!
=====================

Vi har r�tt f� utvecklare vilket tyv�rr inneb�r att arbetet fortskrider r�tt
l�ngsamt. Vi beh�ver helt enkelt mer folk som kan hj�lpa oss! Det finns m�ngder
med uppgifter i behov av dedicerade utvecklare, i alla former fr�n stora projekt
till sm�, fr�n st�d f�r h�rdvara till h�gniv� systemprogrammering och applikationer.
Kort sagt s� finns det n�got f�r alla som kan hj�lpa, oavsett hur duktig du
�r p� programmering.

F�r er som inte �r programmerare s� finns det ocks� m�ngder med saker som ni kan
hj�lpa till med! Bland annat skriva dokumentation, �vers�tta program och dokumentation
till olika spr�k, skapa snygg grafik eller hitta buggar.
Dessa uppgifter �r lika viktiga som programmering!
