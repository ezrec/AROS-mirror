H�r �r Freetype Manager, som anv�nds f�r att installera och konfigurera
nya Truetype-typsnitt i systemet. Inte s� anv�ndarv�nligt, men du kan pilla
p� varje liten detalj. �nnu viktigare, det fungerar. :-)
