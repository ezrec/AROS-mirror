Adam Chodorowski poserar för kameran; iklädd sina hemska
solglasögon som han insisterar att de inte är hans egna. ;-)
