Adam Chodorowski har tagit sig tid att göra ett bra paket av PNG-ikoner, baserade
på Gnome "Gorilla"-ikonpaket, för att visa denna nya AROS-funktion. Du kan även
se det nya "Wanderer preference program", som just nu låter dig ändra bakgrunden
av skrivbordet och mappar i fönster, som även senare kommer tillåta att ändra
alla andra funktioner i Wanderer.

Notera även att alla typsnitt använder antialias.
