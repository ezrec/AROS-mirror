2003-11-24
----------

UAE, Zune och gcc.
