En till bild av Ola utanf�r sitt hem i Norge.
