Mer sidor i Zune-inst�llningar, s� du kan konfigurera anv�ndarinterfacet
precis som *du* vill ha det.
