.. raw:: html

   <table style="text-align: justify; width: 100%;" background="/images/bgcolormain.png" border="0" cellpadding="1" cellspacing="1"><tr><td style="vertical-align: top;">

.. Include:: introduction/index-abstract.sv

`L�s mer... <introduction/index>`__

.. raw:: html

   </td></tr></tbody></table><br>


.. raw:: html

   <table style="width: 100%; text-align: justify; margin-left: auto; margin-right: auto;" background="/images/bgcolormain.png" border="0" cellpadding="1" cellspacing="1"><tr><td>

.. Include:: documentation/developers/contribute-abstract.sv

`L�s mer... <documentation/developers/contribute>`__

.. raw:: html

   </td></tr></table>


.. raw:: html

   <table style="width: 100%; text-align: justify; margin-left: auto; margin-right: auto;" border="0" cellpadding="1" cellspacing="1"><tr><td>

.. Include:: news/index.sv

.. raw:: html

   </td></tr></table><br>


.. raw:: html

   <td style="width: 243px; vertical-align: top;"><table style="text-align: justify; width:100%;" background="/images/bgcolorright.png" border="0" cellpadding="1" cellspacing="1"><tr><td>
   <?php if ($win_ie56) { echo "<img alt=\"Direct download Icon\" src=\"/images/directdownloadicon.gif\" align=\"middle\">";} 
   else { echo "<img alt=\"Direct download Icon\" src=\"/images/directdownloadicon.png\" align=\"middle\">";} ?>Direct Downloads:<br>
   <img style="width: 238px; height: 2px;" alt="spacer" src="images/sidespacer.png"><br>
   Nightly builds skapas automatiskt varje natt, direkt fr�n den senaste k�llkoden. Om du vill prova en AROS live CD, ladda ner "boot ISO" f�r din plattform (i386 or PPC).<br><br>
   <?php virtual("/cgi-bin/files2") ?> <br></td></tr></tbody></table>
   <table style="text-align: justify; width: 100%;" background="/images/bgcolorright.png" border="0" cellpadding="1" cellspacing="1"><tr><td>
   <?php if ($win_ie56) { echo "<img alt=\"Community Icon\" src=\"/images/communityicon.gif\" align=\"middle\">"; } 
   else { echo "<img alt=\"Community Icon\" src=\"/images/communityicon.png\" align=\"middle\">"; } ?> 
   Senaste inl�ggen p� AROS-EXEC forumet:<br><img style="width: 238px; height: 2px;" alt="spacer" src="images/sidespacer.png"><br>
   <a href=http://www.aros-exec.org>AROS-EXEC</a> �r den prim�ra AROS community-sidan. H�r kan du f� hj�lp, h�lla koll p� vad som h�nder inom AROS-v�rlden och posta dina tankar om AROS.<br><br>
   <?php include("/home/groups/a/ar/aros/htdocs/rsfeed/aeforum.php"); ?><br></td></tr></tbody></table>
   <table style="text-align: justify; width: 100%;" background="/images/bgcolorright.png" border="0" cellpadding="1" cellspacing="1"><tr>
   <td style="vertical-align: top;"><?php if ($win_ie56) { echo "<img alt=\"Open Bounty Icon\" src=\"/images/bountyicon1.gif\" align=\"middle\">";} 
   else { echo "<img alt=\"Open Bounty Icon\" src=\"/images/bountyicon1.png\" align=\"middle\">"; } ?>
   �pnna Bounties:<br><img style="width: 177px; height: 2px;" alt="spacer" src="images/sidespacer.png"><br>
   <a href=http://www.teamaros.org>Team AROS</a> �r en supportkampanj f�r AROS som f�rs�ker fungera som en motor f�r AROS-utveckling. Detta g�rs prim�rt genom att samla in donationer f�r specifika projekt.
   <?php include("/home/groups/a/ar/aros/htdocs/rsfeed/teamarosopenb.php"); ?><br></td></tr></table>
   <table style="text-align: justify; width: 100%;" background="/images/bgcolorright.png" border="0" cellpadding="1" cellspacing="1"><tr><td style="vertical-align: top;">
   <?php if ($win_ie56) { echo "<img alt=\"Assigned Bounty Icon\" src=\"/images/bountyicon2.gif\" align=\"middle\">"; } 
   else { echo "<img alt=\"Assigned Bounty Icon\" src=\"/images/bountyicon2.png\" align=\"middle\">"; } ?> 
   Tilldelade Bounties:<br><img style="width: 177px; height: 2px;" alt="spacer" src="images/sidespacer.png"><br>
   <?php include("/home/groups/a/ar/aros/htdocs/rsfeed/teamarosassigned.php"); ?><br></td></tr></table>
   <table style="width: 100%; text-align: justify; margin-left: auto; margin-right: auto;" background="/images/bgcolorright.png" border="0" cellpadding="1" cellspacing="1"><tr><td style="vertical-align: top;">
   <?php if ($win_ie56) { echo "<img alt=\"Syndication Icon\" src=\"/images/rssicon1.gif\" align=\"middle\">"; } else { echo "<img alt=\"Syndication Icon\" src=\"/images/rssicon1.png\" align=\"middle\">"; } ?>
   Syndication Feeds:<br><img style="width: 177px; height: 2px;" alt="spacer" src="images/sidespacer.png"><br>
   <?php  include("/home/groups/a/ar/aros/htdocs/rsfeed/synfeed.php");  ?><br></td></tr></table>
   <table style="text-align: justify; width: 100%;" background="/images/bgcolorright.png" border="0" cellpadding="1" cellspacing="1"><tr><td>
   <?php if ($win_ie56) { echo "<img alt=\"Archive Icon\" src=\"/images/archivedownloadicon.gif\" align=\"middle\">"; } 
   else { echo "<img alt=\"Archive Icon\" src=\"/images/archivedownloadicon.png\" align=\"middle\">"; } ?>
   Latest ARCHIVE submissions:<br><img style="width: 238px; height: 2px;" alt="spacer" src="images/sidespacer.png"><br>
   P� <a href=http://archives.aros-exec.org>The AROS archives</a> hittar du det nyaste materialet f�r AROS, h�r hittar du program, teman, grafik och ytterligare dokumentation.<br><br>
   <?php include("/home/groups/a/ar/aros/htdocs/rsfeed/archives.php"); ?><br></td></tr></table></td></tr></table>
