H�r �r ett fr�nt ritprogram av Hogne "M0ns00n" Titlestad, Lunapaint v0.2.3 (http://www.sub-ether.org/lunapaint) i utveckling. Nu �r tatatype-laddning klart... Mer f�r�ndringar kommer.
