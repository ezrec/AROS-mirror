Adam p� AmiGBG 2002 fair, skrivandes p� sin b�rbara dator.
