===========
Nerladdning
===========

.. Contents::

.. Note::

   N�r du laddar ner "nightly builds", s� m�ste du anv�nda en nerladdnings-
   hanterare s� att du kan �teruppta en avbruten nerladdning, eller en
   textbaserad applikation som t.ex. wget (Du kan anv�nda "wget -c" f�r
   att �teruppta nerladdningen av en fil som �r nerladdad av ett annat program).

Snapshots
=========

Fr�n den 1:a mars 2007 �r snapshots av AROS inte l�ngre tillg�ngliga. Vi
uppmanar alla som vill testa AROS att ladda ner den senaste "nightly build"
ist�llet. AROS v�xer v�ldigt fort, och snapshots inneh�ller oftast
f�r�ldad kod. Vi tror ocks� att "nightly builds" �r mer anv�ndbara med 
tanke p� betatestningen: anv�nd g�rna `bug tracker`__ f�r att rapportera buggar.

__ http://sourceforge.net/tracker/?atid=439463&group_id=43586&func=browse


Nightly builds
==============

"Nightly builds" g�rs, som man ser p� namnet, automatiskt varje natt direkt
fr�n subversions-tr�det och inneh�ller den senaste koden. Men dessa har inte
blivit testade och kan inneh�lla buggar. Dock fungerar dom f�r det mesta bra.

Rapportera g�rna buggar som du hittar n�r du anv�nder "nightly builds" till
`bug tracker`__. F�r �vriga �renden eller fr�gor, kontakta oss via
`AROS-Exec`__ forumen.

.. raw:: html

   <?php virtual( "/cgi-bin/files?type=nightly&lang=sv" ); ?>

__ http://sourceforge.net/tracker/?atid=439463&group_id=43586&func=browse
__ http://aros-exec.org/

