Henning Kiel framf�r logotypen vid entr�n p� IAC (instituto
de Astrofis&iacute;ca de Canarias) i Teneriffa, Spanien.
