Här är ett fränt ritprogram av Hogne "M0ns00n" Titlestad, Lunapaint v0.2.3 (http://www.sub-ether.org/lunapaint) i utveckling. Nu är tatatype-laddning klart... Mer förändringar kommer.
