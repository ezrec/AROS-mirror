Sebastian "Bearly" Heutling som firar sitt arbete med trackdisk.device :).
