V�ntar som m�nga andra p� Amiga Inc p� WoA 1999.
