Fabia Alemagna och Aaron Digulla i cafét 'Dolce Sosta' på ön Ischia
(nära Naples i Italien).
