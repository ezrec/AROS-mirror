2004-03-08
----------

PNG-ikoner och PCI handling tool.
