MesaGL v 6.5 alpha som utvecklas av Kalamatee. Inte så vacker skärmdump, men den senaste dock.
