Tv� instanser av UAS som k�rs samtidigt, som visar b�de Picasso96 och 
chipset-emulation. UAE f�r AROS �r en Zine-applikation, grafik output och 
-input-hanteringen g�rs med hj�lp av en custom class som �r skriven 
just f�r denna hantering.

Ett fullt kvalificerat GUI utvecklas av Adam Chodorowski.
