About(Om) dialogrutan var nyss uppdaterad f�r att visa �nnu mer information,
inte endast f�r att vara extremt h�nf�rande. Du kan �ven se den fina ACSII-logotypen
av Jostein "Taxi" Klemmetsrud som anv�nds nr bilden inte �r tillg�ngligt (Till
exempel p� diskett).
