Adam på AmiGBG 2002 fair, skrivandes på sin bärbara dator.
