H�r visas vinnarna i bakgrundsbildst�vlingen, integrerade i v�ra "nightly builds".
