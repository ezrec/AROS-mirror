==================
Kontaktinformation
==================

:Authors:   Adam Chodorowski, Matthias Rustler 
:Copyright: Copyright � 1995-2009, The AROS Development Team
:Version:   $Revision$
:Date:      $Date$
:Status:    Done.

.. Contents::


Kontakperson
============
Den prim�ra kontaktpersonen f�r teamet som utvecklar AROS �r Aaron "Optimizer"
Digulla. Om du vill ha kontakt med AROS som projekt, till exempel f�r att diskutera
sponsoravtal eller andra former av samarbete, s� �r det personen att kontakta.
Du kan n� honom genom att skicka email till `digulla@aros.org`__.

__ mailto:digulla@aros.org


Mailinglistor
=============

Det finns ett antal AROS-relaterade mailinglistor, vilka �r de viktigaste kanalerna
f�r information och diskussion om AROS f�r utvecklare. F�ljande mailinglistor finns
tillg�ngliga:

+ `AROS Developer`__

  Det h�r �r listan f�r utvecklare d�r diskussioner om utvecklingen av AROS sker.
  H�r postas ocks� statusen fr�n den nattliga kompileringen av AROS. Det �r 
  **starkt** rekommenderat att utvecklare g�r med i den h�r listan eftersom det
  annars �r sv�rt att h�lla sig uppdaterad med den senaste utvecklingen.
  Eftersom det inte finns s� m�nga utvecklare inom AROS, s� �r m�ngden email
  ganska liten men den kan bli ganska h�g om en het diskussion kommer ig�ng.

  .. Note:: Beg�ran om prenumeration p� den h�r listan hanteras inte automatiskt
            utan varje beg�ran kontrolleras av listans administrat�rer. Detta
            inneb�r att det kan ta ett litet tag fr�n det att du skickar in 
            en beg�ran tills dess att du blir en medlem.
  
+ `AROS CVS`__

  P� denna lista f�r utvecklare postas loggar fr�n Subversion-servern s� fort n�got
  s�nder in �ndringar ("commit"). I motsats till den dagliga samlings-loggen som 
  postas p� AROS Developer-listan, d�r varje mail inneh�ller hela dagens aktiviteter
  p� Subversion-servern, s� skickas det separata email f�r varje ins�nd �ndring
  *omedelbart* f�r varje loggad aktivitet. S� om du vill ha n�stan realtids-information
  om vad som h�nder p� Subversion-servern s� �r det h�r listan f�r dig.
  Volymen av mail p� denna lista kan vara ganska h�g.

+ `AROS Website`__

  Skriptsystemet som skapar hemsidan skickar mail till den h�r listan.
  De som jobbar med dokumentationen eller kan laga saker om  n�got h�nder
  med websidan b�r prenumerera p� denna.

F�lj l�nkarna till de administrativa sidorna f�r information om hur man
prenumererar, avbryter prenumerationerer, listarkiv och andra anv�ndbara
funktioner.

__ https://www.hepe.com/mailman/listinfo/aros-dev/
__ http://lists.sourceforge.net/mailman/listinfo/aros-cvs
__ http://lists.sourceforge.net/mailman/listinfo/aros-website

.. _`buggdatabasen`: http://sourceforge.net/tracker/?atid=439463&group_id=43586&func=browse


Forum
=====

AROS-Exec__ �r den officella community-portalen f�r AROS. H�r finner du de
senaste nyheterna om AROS, diskussionsforum, bildgallerier och mycket mer. Det
�r den perfekta m�tesplatsen f�r AROS-anv�ndare fr�n hela v�rlden.

__ http://aros-exec.org/

IRC-Kanaler
===========

Det finns en officiell IRC-kanal f�r AROS, f�ga f�rv�nande d�pt till `#aros`__, p�
FreeNode__-n�tverket. V�nligen anslut till `irc.freenode.net`__ som vidarebefodrar 
dig till en server n�ra dig. Den �r till f�r att diskutera allt m�jligt som �r relaterat
med AROS inklusive utveckling och planer att ta �ver v�rlden. Vid s�llsynta tillf�llen
n�r det �r v�ldigt mycket prat i huvudkanalen flyttar diskussioner relaterade till
utveckling till `#aros.dev`__.

__ irc://irc.freenode.net/aros
__ http://www.freenode.net/
__ irc://irc.freenode.net/
__ irc://irc.freenode.net/aros.dev
