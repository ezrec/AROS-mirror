Fabio Alemagna i sin tr�dg�rd som tar kort mest f�r skoj skull (�ven om han inte verkar tycka
det �r s� kul...) :)
