Fabio Alemagna i sin trädgård som tar kort mest för skoj skull (Även om han inte verkar tycka
det är så kul...) :)
