Här är arbeten av Kalamatee: Konceptionellt GUI för W.I.P AROSTCP Config Tool. Profilsidan låter dig välja/importera/exportera en komplett nätverksprofil/konfiguration. Den tillåter även inställningar i Env-variablerna vilket påverkar AROSTCP.
