Adam Chodorowski poserar f�r kameran; ikl�dd sina hemska
solglas�gon som han insisterar att de inte �r hans egna. ;-)
