Editering i Startup-Sequence med hj�lp av JanoEditor, som f�r tillf�llet
�r AROS standardiserade text-editor.
