Fabia Alemagna och Aaron Digulla i caf�t 'Dolce Sosta' p� �n Ischia
(n�ra Naples i Italien).
