En till bild av Ola utanför sitt hem i Norge.
