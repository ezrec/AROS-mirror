Om du någonsin undrat över hur Fabias ansikte ser ut, så vet du det nu! :)
