Adam Chodorowski har tagit sig tid att g�ra ett bra paket av PNG-ikoner, baserade
p� Gnome "Gorilla"-ikonpaket, f�r att visa denna nya AROS-funktion. Du kan �ven
se det nya "Wanderer preference program", som just nu l�ter dig �ndra bakgrunden
av skrivbordet och mappar i f�nster, som �ven senare kommer till�ta att �ndra
alla andra funktioner i Wanderer.

Notera �ven att alla typsnitt anv�nder antialias.
