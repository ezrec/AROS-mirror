2006-09-01
----------

Här är en del projekt från 2006. AROS visar vårat fräna ritprogram av Hogne "M0ns00n" Titlestad, Lunapaint v0.2.3.  AROS-program har även blivit översatta till ryska. Ett annat projekt av Kalamatee: Konceptiellt GUI för W.I.P AROSTCP Config Tool and MesaGL. Även kommande GUI FTP Client av Suppah (aka voidstar).
