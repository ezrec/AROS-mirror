Henning Kiel framför logotypen vid entrén på IAC (instituto
de Astrofis&iacute;ca de Canarias) i Teneriffa, Spanien.
