Mannen, myten, legenden: nagger (l�s: organizer), evangelist (l�s:
relations-kille) och #AROS IRC channel operator extraordinair�.
