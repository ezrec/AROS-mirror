Tids-inst�llnings-applikationen, klockan och WritePixelArrayAlpha testprogrammen
som visar alpha blending.
