På jobbet.
