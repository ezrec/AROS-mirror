H�r �r arbeten av Kalamatee: Konceptionellt GUI f�r W.I.P AROSTCP Config Tool. Profilsidan l�ter dig v�lja/importera/exportera en komplett n�tverksprofil/konfiguration. Den till�ter �ven inst�llningar i Env-variablerna vilket p�verkar AROSTCP.
