2007-11-30
----------

Under h�sten 2007 har AROS f�tt ett nytt utseende med teman och nya bakgrundsbilder,
ny installer samt att mycket jobb �r gjort inom �vers�ttningar. Mer sk�rmdumpar kommer ...
