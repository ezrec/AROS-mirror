2006-09-01
----------

H�r �r en del projekt fr�n 2006. AROS visar v�rat fr�na ritprogram av Hogne "M0ns00n" Titlestad, Lunapaint v0.2.3.  AROS-program har �ven blivit �versatta till ryska. Ett annat projekt av Kalamatee: Konceptiellt GUI f�r W.I.P AROSTCP Config Tool and MesaGL. �ven kommande GUI FTP Client av Suppah (aka voidstar).
