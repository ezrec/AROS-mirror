Ett f�nster med den nya AROS-installern fr�n Neil Cafferkey.
