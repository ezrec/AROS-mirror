En bunt AROS-utvecklare och AROS-fans, i ett soligt och v�ldigt hett Naples.
