Ett experiment som unders�ker hur m�nga program som du kan trycka in
i en AROS sk�rmdump. Ganska m�nga som du kan se...
