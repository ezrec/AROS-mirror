Tack vare Sergey Mineychev, s� �r alla AROS-programmens cataloger lokaliserade samt att typsnitten �r inlagda (med tillst�nd av Michael Malyshev, ATO).
