==========
Utvecklare
==========

