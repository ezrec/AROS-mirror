MesaGL v 6.5 alpha som utvecklas av Kalamatee. Inte s� vacker sk�rmdump, men den senaste dock.
