====================
AROS p� Amiwest 2012
====================

:F�rfattare:   Jason McMullan
:Datum:        2012-11-02

Vid AmiWest 2012, demonstrerade Samuel Crow and Jason McMullan AROS v1 p� en
Sam460ex fr�n `ACube`__, och FPGA Arcade Replay fr�n `FPGA Arcade`__, samt
Raspberry PI fr�n `Raspberry PI Foundation`__.

Jason McMullan h�ll en ca: 20 minuter l�ng `presentation`__ om ursprunget
till och nuvarande utvecklingsstatus av AROS projektet, och deltog senare
�ven i diskussionspanelen g�llande nul�ge och framtiden f�r Amiga familjens
olika operativsystem.

P� showen delades det �ven ut, DVDs med `Icaros`__ (pc-i386, ABI v0) och
`AROS Vision`__ (amiga-m68k) till alla nya bes�kare.


__ http://acube-systems.biz
__ http://www.fpgaarcade.com
__ http://www.raspberrypi.org

__ http://www.evillabs.net/AROS/AmiWest-2012-Presentation.pdf

__ http://vmwaros.blogspot.com/
__ http://www.natami-news.de/html/aros_vision.html
